module priority_enc_8x3(a,b,v);//{
	input [7:0]a;
	output reg [2:0]b;
	output reg v;

	always @(*) begin//{
		v = 1;
		b = 3'bXXX;
		casex(a)
			8'b00000001 : b = 3'b000;
			8'b0000001x : b = 3'b001;
			8'b000001xx : b = 3'b010;
			8'b00001xxx : b = 3'b011;
			8'b0001xxxx : b = 3'b100;
			8'b001xxxxx : b = 3'b101;
			8'b01xxxxxx : b = 3'b110;
			8'b1xxxxxxx : b = 3'b111;
			default     : v = 0;
		endcase
	end//}
endmodule //}
